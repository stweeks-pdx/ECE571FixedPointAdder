import floatingpointpkg::*;

module FloatingPointAdder(input float AddendA,
			  input float AddendB,
			  input logic Go,
			  output float Result,
			  output logic Zero, 
			  output logic Inf,
			  output logic Nan);
parameter VERSION = "0.1";

endmodule

